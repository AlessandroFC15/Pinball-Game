library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY VGA IS
	PORT(
		CLOCK_24 : IN STD_LOGIC_VECTOR(1 downto 0);
		VGA_HS, VGA_VS : OUT STD_LOGIC;
		VGA_R, VGA_G, VGA_B : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		KEY : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		LED: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END VGA;

ARCHITECTURE MAIN OF VGA IS
	SIGNAL VGACLK, RESET : STD_LOGIC := '0';
	------------------------------------------------------
	COMPONENT PLL1 IS
		PORT(
			CLK_IN_CLK : IN STD_LOGIC := 'X'; -- CLK
			RESET_RESET : IN STD_LOGIC := 'X'; -- RESET
			CLK_OUT_CLK : OUT STD_LOGIC -- CLK
		);
	END COMPONENT PLL1;
	------------------------------------------------------
	COMPONENT SYNC IS
		PORT(
			CLK : IN STD_LOGIC;
			HSYNC, VSYNC : OUT STD_LOGIC;
			R, G, B : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			KEYS : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			LED: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);
	END COMPONENT SYNC;
	
	BEGIN
	
	C1 : SYNC PORT MAP( VGACLK, VGA_HS, VGA_VS, VGA_R, VGA_G, VGA_B, KEY, LED);
	C2 : PLL1 PORT MAP(CLOCK_24(0), RESET, VGACLK);
END MAIN;