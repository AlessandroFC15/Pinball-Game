// PLL1.v

// Generated using ACDS version 13.1 162 at 2017.01.30.16:03:13

`timescale 1 ps / 1 ps
module PLL1 (
		input  wire  clk_in_clk,  //  clk_in.clk
		input  wire  reset_reset, //   reset.reset
		output wire  clk_out_clk  // clk_out.clk
	);

	PLL1_altpll_0 altpll_0 (
		.clk       (clk_in_clk),  //       inclk_interface.clk
		.reset     (reset_reset), // inclk_interface_reset.reset
		.read      (),            //             pll_slave.read
		.write     (),            //                      .write
		.address   (),            //                      .address
		.readdata  (),            //                      .readdata
		.writedata (),            //                      .writedata
		.c0        (clk_out_clk), //                    c0.clk
		.areset    (),            //        areset_conduit.export
		.locked    (),            //        locked_conduit.export
		.phasedone ()             //     phasedone_conduit.export
	);

endmodule
